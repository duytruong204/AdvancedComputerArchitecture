`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/00_mux/mux_2to1_1bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/00_mux/mux_2to1_2bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/00_mux/mux_2to1_3bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/00_mux/mux_2to1_4bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/00_mux/mux_2to1_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/00_mux/mux_4to1_1bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/00_mux/mux_4to1_4bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/00_mux/mux_4to1_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/00_mux/mux_8to1_1bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/00_mux/mux_8to1_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/00_mux/mux_16to1_1bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/00_mux/mux_16to1_32bit.sv"

`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/01_operation/full_adder_1bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/01_operation/full_adder_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/01_operation/sll_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/01_operation/slt_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/01_operation/sltu_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/01_operation/sra_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/01_operation/srl_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/01_operation/xor_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/01_operation/or_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/01_operation/and_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/01_operation/equal_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/01_operation/equal_20bit.sv"

`include "D:/Application/altera/13.0sp1/Project/Single_Cycle_RISC_V/milestone2_ver1/00_src/00_common/02_memory/memory.sv"