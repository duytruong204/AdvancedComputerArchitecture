// Mux
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_2to1_1bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_2to1_2bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_2to1_3bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_2to1_4bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_2to1_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_2to1_nbit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_4to1_1bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_4to1_2bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_4to1_4bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_4to1_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_8to1_1bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_8to1_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_16to1_1bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/00_mux/mux_16to1_32bit.sv"
// operation
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/full_adder_1bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/full_adder_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/full_adder_nbit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/sll_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/slt_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/sltu_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/sra_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/srl_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/xor_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/or_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/and_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/equal_32bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/equal_20bit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/01_operation/equal_nbit.sv"
// memory
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/02_memory/d_flip_flop.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/02_memory/memory.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/02_memory/single_port_ram.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/00_common/02_memory/memory_ram.sv"
// sub block
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/01_sub_block/alu.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/01_sub_block/brc.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/01_sub_block/control_logic.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/01_sub_block/imm_gen.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/01_sub_block/inst_mem.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/01_sub_block/lsu.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/01_sub_block/pc.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/01_sub_block/regfile.sv"
// pipeline registers
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/02_pipelined_regs/IF_ID_reg.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/02_pipelined_regs/ID_EX_reg.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/02_pipelined_regs/EX_MEM_reg.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/02_pipelined_regs/MEM_WB_reg.sv"
// pipelined control
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/03_pipelined_control/branch_taken.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/03_pipelined_control/stall_flush_unit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/03_pipelined_control/load_pending.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/03_pipelined_control/forwarding_unit.sv"
`include "D:/Application/altera/13.0sp1/Project/Pipeline_RISC_V/pipelined_branch_prediction/00_src/03_pipelined_control/branch_prediction_unit.sv"